module writeback(
    input [3:0] icode,      
    input [3:0] valA,        
    input [3:0] valB,
    input [63:0] valE,          
    input [63:0] valP,
    input [63:0] valM,
    
);

endmodule